--Τύποι που ορίζονται από τον χρήστη (user-defined types)
--Εκτός από τους προκαθορισμένους και προτυποποιημένους τύπους δεδομένων που
--ο κάθε χρήστης μπορεί να δημιουργήσει τους δικούς του τύπους
--δεδομένων, ώστε να χειριστεί πιο εύκολα τη σχεδίαση ενός συστήμαος. Η δήλωση του τύπου
--δεδομένων μπορεί να γίνει στο σώμα δηλώσεων της αρχιτεκτονικής ή σε ξεχωριστό πακέτο
--(package), όπως είναι και το πιο βολικό σε μεγάλες σχεδιάσεις. Η δήλωση ενός τύπου δεδομένων
--από το χρήστη γίνεται με την εξής γενική μορφή:
TYPE όνομα_τύπου IS περιγραφή τύπου;

--Ακέραιοι τύποι ορισμένοι από τον χρήστη
--συγκεκριμένο σύνολο ακέραιων τιμών
TYPE όνομα_τύπου IS RANGE αρχική_τιμή ΤΟ τελική_τιμή;

Παράδειγμα:
TYPE temperature IS RANGE 0 TO 273;
SIGNAL s : temperature;
