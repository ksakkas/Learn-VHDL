ENTITY full_adder IS 
PORT (cin, a, b : IN BIT; 
		s, cout : OUT BIT); 
END full_adder;
