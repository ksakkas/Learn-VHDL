--Τύποι standard logic (πακέτο std_logic_1164)

--Όλες οι τιμές που λαμβάνει ένα σήμα std_logic είναι οι εξής:
-- '0' Λογικό μηδέν
-- '1' Λογικό ένα
-- 'Ζ' Υψηλή εμπέδηση
-- '-' Αδιάφορη κατάσταση
-- 'U' Μη αρχικοποιημένη κατάσταση (Uninitialized)
-- 'X' Άγνωστη κατάσταση
-- 'L' Ασθενής χαμηλή (Weak low)
-- 'H' Ασθενής υψηλή (Weak high)
-- 'W' Ασθενής άγνωστη (Weak unknown)