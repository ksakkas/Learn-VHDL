--Υποτύποι δεδομένων
--Οι υποτύποι ορίζουν μια ειδική υποκατηγορία ενός τύπου δεδομένων. Για παράδειγμα, μπορούμε
--να ορίσουμε ως υποτύπο του τύπου SIGNED, αυτόν που περιγράφει σήματα που λαμβάνουν
--προσημασμένες τιμές με οκτώ bits:

SUBTYPE sample IS SIGNED(7 downto 0);

SIGNAL normal : sample;