--Ο απαριθµητής είναι ένα ακουθιακό κύκλωµα, που αυξάνει την
--έξοδό του κατά ένα κάθε φορά που δέχεται ένα παλµό ρολογιού. Για το συγχρονισµό
--διεργασιών µε µεταβάσεις σηµάτων (όπως ο παλµός clock) η γλώσσα VHDL χρησιµοποιεί µια
--δοµή που ονοµάζεται PROCESS (διεργασία). Οι εντολές που περιλαµβάνονται στην PROCESS,
--όπως για παράδειγµα η IF, εκτελούνται σειριακά, αλλά οι αναθέσεις των σηµάτων
--γίνονται µόνον στο τέλος, µε σύγχρονο τρόπο. 

LIBRARY ieee;                        --Δήλωση Βιβλιοθήκης
USE ieee.std_logic_1164.all;         --Δήλωση πακέτων
USE ieee.std_logic_unsigned.all;     --Δήλωση πακέτων


-----------------------------------------------------------------------------------------


ENTITY counter IS                    --Δήλωση οντότητας με όνομα counter
--Η δήλωση των διασυνδέσεων γίνεται µε τη βοήθεια της κωδικής δήλωσης PORT (…), όπου
--µέσα στην παρένθεση γίνονται οι δηλώσεις των σηµάτων διασύνδεσης:
--• ΙΝ Χρησιµοποιείται για σήµατα που αποτελούν εισόδους στη βαθµίδα
PORT(clk : IN std_logic;             --Δήλωση clk ως ακέραια 
--Όπως φαίνεται στο µέρος της οντότητας, ο
--απαριθµητής έχει είσοδο παλµών ρολογιού (clk). H είσοδος αυτή είναι σήµα του τύπου
--std_logic, που όπως θα δούµε ορίζει ένα σύνολο εννέα τιµών, τις οποίες µπορεί να λάβει ένα
--σήµα. Οι κυριότερες είναι οι '1', '0', 'Ζ', που η κάθε µια ορίζεται ως ένας χαρακτήρας. 
q : OUT std_logic_vector (3 DOWNTO 0));
--Η έξοδος q ορίζεται ως ένα σήµα τύπου std_logic_vector, δηλαδή ως ένας πίνακας
--χαρακτήρων τύπου std_logic. Το (3 downto 0) στη δήλωση του τύπου σηµαίνει ότι το
--σήµα έχει 4 bit. Τα στοιχεία του πίνακα είναι τα q(3), q(2), q(1), q(0), µε πρώτο εξ’
--αριστερών το πιο σηµαντικό bit
END counter;                       --Τέλος οντότητας


----------------------------------------------------------------------------------------


ARCHITECTURE behaviour OF counter IS        --Δήλωση αρχιτεκτονικής με όνομα behaviour απο την οντότητα counter
SIGNAL m : std_logic_vector (3 DOWNTO 0);   --Δήλωση σήματος με όνομα m τύπου vector (μεγάθους 4) 
BEGIN                                       --Αρχή
PROCESS(clk)                                --Διεργασία clk
BEGIN                                       --Αρχή
IF clk 'event AND clk='1' THEN              --Αν το clk έχει παλμό και είναι 1 (άνοδος) τότε
m<= m+1;                                    -- m = m + 1
ELSE                                        --Αλλιώς
m<=m;                                       --m = m
END IF;                                     --Τέλος if
END process;                                --Τέλος διεργασίας
q<=m;                                       --q = m
END behaviour;                              --Τέλος αρχιτεκτονικής