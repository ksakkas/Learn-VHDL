--Τελεστές ανάθεσης
-- <=    Αναθέτει τιμές σε σήματα    <όνομα_σήματος> <= <έκφραση>     s1<=s2+s3;
-- :=    Αναθέτει τιμές σε μεταβλητές (δίνει αρχικές τιμές σε σήματα, κατά τη δήλωσή τους)
--       <όνομα_μεταβλητής> :=<έκφραση>     v1 := s1 OR s2;     v2 := "1010";
-- =>    Δίνει τιμές σε στοιχεία πινάκων   v3:=(0=>'1', 1=>'0', OTHERS=>'0');

--Λογικοί τελεστές
--Not Αντιστροφή
--And Και
--Nand Όχι Και
--Or Ή
--Nor Ούτε
--Xor Αποκλειστικό Ή
--Xnor Αποκλειστικό Ούτε

--Σχεσιακοί τελεστές
-- = Ισότητα
-- /= (ιάφορο
-- < Μικρότερο
-- <= Μικρότερο ή ίσο
-- > Μεγαλύτερο
-- >= Μεγαλύτερο ή ίσο