--H εντολή SELECT
--Μια βασική σύγχρονη εντολή είναι η SELECT, που συντάσσεται ως εξής:
WITH αναγνωριστικό SELECT
Έκφραση_ανάθεσης_τιμής WHEN τιμή
Ανάθεση_τιμής WHEN τιμή
Ανάθεση_τιμής WHEN τιμή
....;

--Το «αναγνωριστικό» μπορεί να είναι το όνομα ενός σήματος. Επειδή η εντολή SELECT
--απαιτεί να καλύπτονται όλες οι δυνατές τιμές που λαμβάνει το «αναγνωριστικό», συχνά η
--παραπάνω δομή κώδικα κλείνει με την έκφραση WHEN OTHERS; στην οποία περιλαμβάνονται
--όλες οι δυνατές τιμές του αναγνωριστικού που δεν έχουν αναφερθεί παραπάνω. Η εντολή
--SELECT προφανώς υλοποιεί κυκλώματα με εισόδους επιλογής, όπως οι πολυπλέκτες, οι
--αποκωδικοποιητές και οι κωδικοποιητές.

--Να σχεδιαστεί πολυπλέκτης δύο καναλιών, όπου το κάθε κανάλι έχει εύρος 8-bit.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
---------------------------------------------------------
ENTITY part2 IS
PORT (Α, Β : IN std_logic_vector (7 downto 0);
s : IN std_logic;
F : OUT std_logic_vector(7 downto 0));
END part2;
----------------------------------------------------------
ARCHITECTURE behaviour OF part2 IS
BEGIN
WITH s SELECT
F<= A WHEN '0',
B WHEN OTHERS;
END behaviour;