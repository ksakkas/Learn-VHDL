--Εντολή LOOP
--Η εντολή LOOP δημιουργεί βρόχους επανάληψης, όπου υλοποιούνται πολλά στιγμιότυπα
--(instances) ενός κυκλώματος. Έτσι, για παράδειγμα, με μια LOOP μπορούμε να επαναλάβουμε
--ένα D Flip-Flop όσες φορές χρειάζεται για τη δημιουργία ενός καταχωρητή. Σε έναν απαριθμητή
--η Loop μπορεί να χρησιμοποιηθεί για την παραγωγή των διαδοχικών αυξήσεων της εξόδου, μέχρι
--να συμπληρωθεί ο απαραίτητος αριθμός καταστάσεων. Σε όλες τις περιπτώσεις, η LOOP πρέπει
--να βρίσκεται μέσα σε διεργασία ή υποπρόγραμμα. Η αντίστοιχη σύγχρονη εντολή είναι η
--GENERATE. Οι μορφές με τις οποίες συναντούμε τη LOOP είναι οι εξής:

--Α. LOOP χωρίς συνθήκη (infinite loop-ατέρμων βρόχος):
[ετικέτα_βρόχου:] LOOP
ακολουθιακός κώδικας
END LOOP [ετικέτα_βρόχου];

--Μοντελοποίηση απαριθμητή mod 16 με εντολή LOOP.
--Ο παρακάτω κώδικας εισάγει έναν ατέρμονα βρόχο LOOP μέσα σε μια διεργασία, με σκοπό την
--αύξηση της εξόδου σε κάθε θετικό μέτωπο ρολογιού, ξεκινώντας από την τιμή μηδέν. Η
--επανάληψη διακόπτεται κάθε φορά στην αρχή, αναμένοντας την εκπλήρωση της συνθήκης
--WAIT. Στο θετικό μέτωπο του σήματος clk η LOOP συνεχίζει, οπότε ανανεώνει την τιμή της
--μεταβλητής m και την έξοδο q. Ας προσεχθεί ό μηδενισμός της m μόλις αυτή αυξηθεί και γίνει
--16. Αυτό πετυχαίνεται με το υπόλοιπο της διαίρεσης (mod) με το 16, που γίνεται μηδέν μονον
--όταν m=16. Τέλος, η διεργασία προφανώς δεν έχει λίστα ευαισθησίας, αφού περιέχεται εντολή
--WAIT.
--Κάθε φορά που αναστέλλεται η διεργασία εξαιτίας της εντολής WAIT, αποδίδονται και οι
--τιμές των σημάτων. Ο παρακάτω κώδικας μοντελοποιεί τη λειτουργία του απαριθμητή, αλλά δεν
--παρέχει κάποιο μηχανισμό για την έξοδο από τον ατέρμονα βρόχο.

------------------------------------
ENTITY loop_counter IS
PORT(clk : IN bit;
q : OUT natural);
END loop_counter;
------------------------------------
ARCHITECTURE behaviour OF loop_counter IS
BEGIN
PROCESS
VARIABLE m : natural :=0;
BEGIN
q<=m;
LOOP
wait until clk'event AND clk ='1';
m:=(m+1) mod 16;
q<=(m);
END LOOP;
END PROCESS;
END behaviour;

--B. LOOP με εντολή EXIT
--Η exit διακόπτει την εκτέλεση του βρόχου και μεταφέρει τη σειρά εκτέλεσης των εντολών έξω
--από το βρόχο. Μπορεί να διατυπωθεί απλά, χωρίς συνθήκη (unconditional) ή με συνθήκη. Η
--γενική διατύπωση έχει ως εξής:
[ετικέτα:] exit [ετικέτα_βρόχου] [when συνθήκη]
--Ως γνωστό, οι αγγύλες σημαίνουν προαιρετική σύνταξη. Ένα γενικό παράδειγμα διατύπωσης
--είναι το εξής:

PROCESS
VARIABLE m : natural;
BEGIN
LOOP
m:=m+1;
exit when m>10;
END LOOP;
--O έλεγχος της εκτέλεσης μεταφέρεται σ’ αυτό το σημείο,
--όταν η συνθήκη m>10 γίνει αληθής
END PROCESS;

--Γ. LOOP με FOR
--Πρόκειται για την πιο διαδεδομένη χρήση της LOOP. Η σύνταξη της εντολής είναι ως εξής:
[ετικέτα:] FOR αναγνωριστικό IN περιοχή_τιμών LOOP
ακολουθιακός κώδικας
END LOOP [ετικέτα];

--Δ. LOOP με WHILE
--H εντολή αυτή συντάσσεται ως εξής:
[ετικέτα:] WHILE συνθήκη LOOP
ακολουθιακός κώδικας
END LOOP [ετικέτα];