--Καταχωρητές
--Ως καταχωρητές θεωρούμε
--ένα σύνολο από Flip Flops, τα οποία είναι κατάλληλα συνδεδεμένα μεταξύ τους και δέχονται ένα
--κοινό ωρολογιακό σήμα. Σε κάθε Flip Flop μπορεί να αποθηκευτεί 1 bit πληροφορίας. Έτσι, σ’
--έναν καταχωρητή ο οποίος αποτελείται από n Flip Flops μπορούμε να αποθηκευτούν n bits
--πληροφορίας. Άρα, για την δημιουργία ενός καταχωρητή χωρητικότητας 8 bits θα πρέπει να
--χρησιμοποιηθούν οκτώ Flip-Flops.

--οι καταχωρητές
--χωρίζονται στις εξής τέσσερις κατηγορίες:
--• Καταχωρητές σειριακής εισόδου-σειριακής εξόδου
--• Καταχωρητές σειριακής εισόδου-παράλληλης εξόδου
--• Καταχωρητές παράλληλης εισόδου-σειριακής εξόδου
--• Καταχωρητές παράλληλης εισόδου-παράλληλης εξόδου

--Να σχεδιαστεί ένας καταχωρητής παράλληλης εισόδου - παράλληλης εξόδου με
--ασύγχρονη είσοδο clear. Ο καταχωρητής να σχεδιαστεί με δήλωση γενικής σταθερής
--(GENERIC) ώστε να μπορεί να επεκταθεί σε οποιοδήποτε εύρος bits.
--Η επέκταση του καταχωρητή σε οποιοδήποτε εύρος bits γίνεται μεταβάλλοντας τον αριθμό των Flip-Flops.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
---------------------------------------------
ENTITY reg IS
GENERIC(N : NATURAL :=8);
PORT (d: IN std_logic_vector(N-1 DOWNTO 0);
clock, clear: IN std_logic;
q: OUT std_logic_vector(N-1 DOWNTO 0));
END reg;
---------------------------------------------
ARCHITECTURE behaviour OF reg IS
BEGIN
PROCESS (clear, clock)
BEGIN
IF clear='0' THEN
q<=(OTHERS=>'0');
ELSIF clock'event AND clock='1' THEN
q<=d;
END IF;
END process;
END behaviour;
