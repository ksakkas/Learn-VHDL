--Απαριθμητές
--Απαριθμητές ονομάζονται τα
--κυκλώματα που μπορούν να αυξήσουν ή να μειώσουν την τιμή της εξόδου τους κατά ένα, όταν
--στην είσοδο ρολογιού δέχονται παλμό clock. Τα κυκλώματα των απαριθμητών μπορούν να
--χρησιμοποιηθούν α) για να μετρούν πόσες φορές εμφανίστηκε κάποιο γεγονός, για παράδειγμα
--πόσες φορές ένα περιφερειακό διακόπτει τον επεξεργαστή β) για την απαρίθμηση διαδοχικών
--εργασιών σε ένα σύστημα, όπως για παράδειγμα για την απαρίθμηση και τον έλεγχο των φάσεων
--εκτέλεσης εντολής σε μικροεπεξεργαστή γ) για την παραγωγή χρονικών καθυστερήσεων, όπως
--σε κυκλώματα χρονιστών.

--Γενικός απαριθμητής με είσοδο παράλληλης φόρτωσης, είσοδο μηδενισμού και
--είσοδο enable.
--Ο απαριθμητής που θα σχεδιάσουμε εδώ, λειτουργεί καταμετρώντας προς τα πάνω (up counter).
--Είναι σχεδιασμένος ως γενικός απαριθμητής mod N, με τη βοήθεια της δήλωσης GENERIC. Για
--Ν=4 ο απαριθμητής λειτουργεί με 4 bits. (ιαθέτει είσοδο μηδενισμού (Resetn) και είσοδο
--ενεργοποίησης (en). Επίσης, διαθέτει είσοδο παράλληλης φόρτωσης Α και ακροδέκτη για την
--ενεργοποίηση της παράλληλης φόρτωσης Ld.
--Όταν N=4, η έξοδος έχει εύρος 4 bits σημαίνει ότι μπορεί να πάρει μέχρι και την τιμή
--“1111”, που στο δεκαδικό σύστημα είναι ο αριθμός 15. (ηλαδή καταμετρά συνολικά δεκαέξι
--καταστάσεις.
--Οι είσοδοι resetn και en είναι οι είσοδοι μηδενισμού και ενεργοποίησης. Εάν η είσοδος
--resetn βρίσκεται σε λογική κατάσταση μηδέν, η έξοδος του κυκλώματος (q) θα μηδενίζεται.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
---------------------------------------------------------------
ENTITY counter IS
GENERIC(N : NATURAL :=8);
PORT(clk, ld, resetn, en : IN std_logic;
A: IN std_logic_vector (N-1 DOWNTO 0);
q: OUT std_logic_vector (N-1 DOWNTO 0));
END counter;
---------------------------------------------------------------
ARCHITECTURE behaviour OF counter IS
SIGNAL m : std_logic_vector (3 DOWNTO 0);
BEGIN
PROCESS(clk, resetn)
BEGIN
IF resent='0' THEN
m<=(OTHERS=>'0');
ELSIF clk'event AND clk='1' THEN
IF en='1' THEN
IF ld='1' THEN
m<=A;
ELSE
m<= m+1;
END IF;
ELSE
m<=m;
END IF;
END IF;
END process;
q<=m;
END behaviour;