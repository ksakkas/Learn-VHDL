library: ieee
