--Η οντότητα (entity) περιγράφει το κύκλωµα ως βαθµίδα, µε εισόδους και εξόδους.
--Περιλαµβάνει µόνο τις διασυνδέσεις που έχει το κύκλωµα µε άλλες βαθµίδες αλλά αποκρύπτει τη
--λειτουργία του κυκλώµατος. Το αναγνωριστικό όνοµα που δίνει ο σχεδιαστής στην οντότητα
--καθώς και τα σήµατα εισόδου και εξόδου είναι καθοριστικά για κάθε υλοποίηση τoυ κυκλώµατος αυτού. 

-- Μετά την κωδική λέξη ENTITY ακολουθεί το όνοµα της οντότητας, 
--που µπορεί να είναι οποιαδήποτε µηδεσµευµένη λέξη και η κωδική λέξη IS:

ENTITY όνοµα_οντότητας IS; 

--Η δήλωση των διασυνδέσεων γίνεται µε τη βοήθεια της κωδικής δήλωσης PORT (…), όπου
--µέσα στην παρένθεση γίνονται οι δηλώσεις των σηµάτων διασύνδεσης: 

PORT(όνοµα_σήµατος_1 : τρόπος_λειτουργίας τύπος_σήµατος_1;
 όνοµα_σήµατος_2 : τρόπος_λειτουργίας τύπος_σήµατος_2;
 ...
 όνοµα_σήµατος_N : τρόπος_λειτουργίας τύπος_σήµατος_N);

 --Ο «τρόπος_λειτουργίας» (mode) καθορίζει την κατεύθυνση του σήµατος διασύνδεσης και
--µπορεί να ανήκει σε µια από τις παρακάτω κατηγορίες:
--• ΙΝ Χρησιµοποιείται για σήµατα που αποτελούν εισόδους στη βαθµίδα
--• OUT Χρησιµοποιείται για σήµατα που αποτελούν εξόδους. Η κατάσταση τέτοιων
--σηµάτων µπορεί να αναγνωριστεί µόνον από άλλες βαθµίδες τις οποίες τα σήµατα
--τροφοδοτούν, όχι όµως από το εσωτερικό της οντότητας
--• INOUT Πρόκειται για δικατευθυντήρια σήµατα, όπως αυτά που συνδέονται µε
--διαδρόµους δεδοµένων δύο κατευθύνσεων (π.χ. σήµατα εισόδου/εξόδου σε µνήµη)
--• BUFFER για σήµατα εξόδου, που ταυτόχρονα µπορούν να διαβαστούν στο εσωτερικό της οντότητας

--Η δήλωση της οντότητας κλείνει µε την πρόταση τέλους:

END [ENTITY] [όνοµα_οντότητας]; 

