--Η γλώσσα VHDL διαχειρίζεται τρία «αντικείμενα δεδομένων» (data objects) τα οποία μπορούν
--να μεταφέρουν πληροφορία μέσα στο σύστημα και να αποδίδουν τιμές σε διάφορα σημεία. Σε
--κάθε αντικείμενο δίνουμε ένα όνομα και το oρίζουμε σύμφωνα με κάποιο «τύπο δεδομένων»
--(data type). Επίσης, κάθε αντικείμενο έχει σε κάθε στιγμή κάποια τιμή. Τα αντικείμενα
--δεδομένων που χρησιμοποιούνται είναι:
--Α. Σήματα (SIGNALS)
--B. Μεταβλητές (VARIABLES)
--Γ. Σταθερές (CONSTANTS)

--Τα σήματα είναι τα πλέον σημαντικά, καθώς αποδίδουν τιμές στα καλώδια του κυκλώματος
--και αντιπροσωπεύουν τις διασυνδέσεις ανάμεσα σε μονάδες του κυκλώματος. Μπορούν να
--χρησιμοποιηθούν τόσο σε τμήματα κώδικα που περιλαμβάνουν σύγχρονες εντολές, όσο και σε
--ακολουθιακά τμήματα κώδικα.

--Οι μεταβλητές χρησιμοποιούνται για την προσωρινή αποθήκευση τιμών που προκύπτουν
--από την τέλεση αριθμητικών πράξεων. Μια μεταβλητή δηλώνεται και χρησιμοποιείται μόνο σε
--τμήματα του κώδικα που περιλαμβάνουν «ακολουθιακές εντολές». Ένα τέτοιο τμήμα κώδικα
--δηλώνεται συνήθως ως ΔΙΕΡΓΑΣΙΑ (PROCESS) και χρησιμοποιείται κυρίως για την περιγραφή
--ακολουθιακών κυκλωμάτων

--Οι σταθερές λαμβάνουν τιμή κατά τη δήλωσή τους και η τιμή αυτή παραμένει στη
--συνέχεια σταθερή. Άρα, η σταθερά δεν αντιπροσωπεύει κάποιο καλώδιο του συστήματος, απλά
--μεταφέρει μια συγκεκριμένη αριθμητική τιμή, όπου χρειάζεται.

