--Η εντολή IF
--Η εντολή Αν είναι εντολή διακλάδωσης υπό συνθήκη. Μπορεί να γραφεί μόνον μέσα σε
--ακολουθιακό τμήμα κώδικα (συνήθως διεργασία-PROCESS). Ελέγχει αν μια συνθήκη είναι
--αληθής, οπότε εκτελεί το μέρος του κώδικα που ακολουθεί, αλλιώς ελέγχει μια νέα σειρά
--συνθηκών και εκτελεί το αντίστοιχο μέρος του κώδικα. Η πλήρης περιγραφή της IF έχει ως
--εξής:
IF συνθήκη THEN
Προτάσεις ανάθεσης;
ELSIF συνθήκη THEN
Προτάσεις ανάθεσης
ELSE
Προτάσεις ανάθεσης;
END IF;

