--Δομικά στοιχεία (components)
--Τα υποκυκλώματα που συμπεριλαμβάνονται σε μια ανώτερη οντότητα (top-level entity)
--ονομάζονται δομικά στοιχεία (components). Τα στοιχεία είναι μικρότερα κυκλώματα, που έχουν
--ήδη περιγραφεί σε VHDL. Τέτοια αρχεία μπορεί να είναι έτοιμοι κώδικες που περιλαμβάνονται
--στο λογισμικό σχεδίασης ή κώδικες που σχεδιάζει ο ίδιος ο χρήστης.
--Τα κύρια χαρακτηριστικά της σχεδίασης μιας ανώτερης ιεραρχικής οντότητας με
--υποκυκλώματα είναι η δήλωση των δομικών στοιχείων που περιέχονται στο κύκλωμα, καθώς και
--η περιγραφή του τρόπου με τον οποίο τα στοιχεία συνδέονται μεταξύ τους.
--Με την δήλωση του κάθε υποκυκλώματος καθορίζουμε το όνομα του, καθώς και τα ονόματα
--των εισόδων και των εξόδων του. Η δήλωση των δομικών στοιχείων μπορεί να γίνει στην
--περιοχή δηλώσεων της αρχιτεκτονικής ή σ’ ένα πακέτο (PACKAGE). Η γενική μορφή μιας
--τέτοιας δήλωσηςείναι ως εξής:
COMPONENT όνομα συνιστώσας
[GENERIC (όνομα παραμέτρου : integer := τιμή; ]
PORT (όνομα ακροδέκτη : mode τύπος;
όνομα ακροδέκτη : mode τύπος );
END COMPONENT;

--Παρακάτω δίνεται ένα παράδειγμα δήλωσης ενός απαριθμητή (οντότητα upcount) ως δομικού στοιχείου:
COMPONENT upcount
PORT(clock, Resetn, E: IN std_logic;
Q: OUT std_logic_vector (3 DOWNTO 0));
END COMPONENT;

--Στη συνέχεια, στο κύριο σώμα της αρχιτεκτονικής, πρέπει να δημιουργήσουμε στιγμιότυπα για
--τα υποκυκλώματα που έχουμε δηλώσει, και να περιγράψουμε τις συνδέσεις τους. Η δημιουργία
--των στιγμιοτύπων γίνεται πάντα μετά τη δήλωση ενός δομικού στοιχείου. Τα στιγμιότυπα είναι της μορφής:
Όνομα_στιγμιότυπου: όνομα στοιχείου PORT MAP (ονόματα σημάτων);
--Στη δήλωση PORT MAP δημιουργούμε τις διασυνδέσεις ανάμεσα στις εισόδους/εξόδους
--κάθε υποκυκλώματος και στα σήματα της ανώτερης οντότητας την οποία περιγράφουμε.
--Η ετικέτα «όνομα_στιγμιότυπου» είναι υποχρεωτική. Η ονομασία μπορεί να είναι
--οποιαδήποτε, αρκεί να υπακούει στους κανόνες ονοματοδοσίας των αναγνωριστικών.

stage1: upcount PORT MAP (clk, Rstn, En, QS);
