entity nor_gate is
port (a , b : in bit;
		y   : out bit);  
end nor_gate;
