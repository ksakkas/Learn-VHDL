--Η εντολή FOR…GENERATE
--Η σύγχρονη εντολή GENERATE δημιουργεί έναν βρόχο όπου επαναλαμβάνεται ένα τμήμα
--κώδικα, με τη βοήθεια ενός δείκτη. Ο κώδικας μπορεί να περιλαμβάνει απλές αναθέσεις
--σημάτων, αριθμητικές πράξεις ή και στιγμιότυπα κυκλωμάτων. Αποτελεί, λοιπόν, ένα δυναμικό
--τρόπο δημιουργίας μεγαλύτερων κυκλωμάτων από απλούστερα και βοηθά στη γραφή
--συμπυκνωμένου κώδικα. Η εντολή GENERATE εμφανίζεται με δύο τρόπους. Ο ένας είναι υπό
--συνθήκη (IF…GENERATE) και ο άλλος χωρίς συνθήκη (FOR…GENERATE). Θα εξεταστεί
--δεύτερος τρόπος, που είναι ο πλέον συνηθισμένος. Η διατύπωση της εντολής είναι ως εξής:

Ετικέτα: FOR αναγνωριστικό ΙΝ περιοχή τιμών GENERATE
Τμήμα σύγχρονων εντολών
END GENERATE;

--Στην παραπάνω διατύπωση, η ετικέτα είναι υποχρεωτική.
--Για παράδειγμα, το παρακάτω τμήμα κώδικα αντιστρέφει τη σειρά των bits σε ένα σήμα x με
--εύρος οκτώ bits και αναθέτει την τιμή σε ένα σήμα y.

SIGNAL x,y,z : std_logic_vector(7 downto 0);
-----------------------------------------
My_label: FOR i IN 0 TO 7 GENERATE
y(i)<=x(7-i);
END GENERATE;

