--Τύποι πινάκων
--Ένας πίνακας μπορεί να είναι μονοδιάστατος ή περισσότερων διαστάσεων και δηλώνεται γενικά
--ως εξής:
TYPE όνομα_τύπου IS ARRAY (περιοχή δεικτών) OF τύπος_στοιχείων;

--Για παράδειγμα ένας πίνακας ακεραίων με πέντε στοιχεία μπορεί να οριστεί ως εξής:
TYPE int_matrix IS ARRAY(1 TO 5) OF INTEGER;

--Μια σταθερά (constant) αυτού του τύπου θα οριστεί ως εξής:
CONSTANT c1: int_matrix(1 TO 5) :=(8, -2, 10, -20, 15);  --c1(1)=8, c1(2)=-2

--Προκειμένου να αφήσουμε ελεύθερη την περιοχή δεικτών να καταλάβει όλο το εύρος των
--ακεραίων από 0 έως το άνω όριο, γράφουμε τη δήλωση:
TYPE my_type IS ARRAY(NATURAL RANGE <>) OF INTEGER;
