--Κάποιοι βασικοί τύποι δεδομένων ανήκουν στην αρχική προτυποποίηση της γλώσσας (πακέτο
--standard της βιβλιοθήκης std) και λειτουργούν χωρίς να χρειάζεται αναφορά σε βιβλιοθήκες.
--Οι βασικοί αυτοί τύποι είναι οι εξής:

--BIT Τα σήματα αυτού του τύπου μπορούν να πάρουν τις τιμές ‘0’ ή ‘1’. Ο τύπος αυτός
--υποστηρίζει λογικούς και σχεσιακούς τελεστές. Θεωρείται βαθμωτός (scalar) τύπος, καθώς
--αποτελείται από ένα bit. Παράδειγμα δήλωσης σήματος τύπου bit:
signal flag : bit;

--BIT_VECTOR Τα σήματα μπορούν να λάβουν μια σειρά τιμών ‘0’ ή ‘1’. (δηλαδή, ο τύπος
--ορίζεται ως ένας μονοδιάστατος πίνακας (array) με στοιχεία BIT. H αλληλουχία των bits
--“10101100” αποτελεί ένα διάνυσμα (vector) με οκτώ στοιχεία. Ο τύπος bit_vector
--υποστηρίζει λογικούς και σχεσιακούς τελεστές, καθώς και τελεστές ολίσθησης και συνένωσης.
--Ένας τρόπος με τον οποίο ορίζεται σήμα αυτού του τύπου δίνεται στο παράδειγμα:
signal data_bus : bit_vector (7 downto 0);

--INTEGER Ένα σήμα αυτού του τύπου μεταφέρει ακέραιες τιμές. Από τη σκοπιά του χρήστη
--είναι βαθμωτός τύπος, καθώς διαχειρίζεται μία μόνο τιμή. Από την άλλη μεριά, σε επίπεδο
--σήματος περιλαμβάνει ένα σύνολο bits. Γενικά, έχει μήκος 32 bits και εύρος τιμών από –(2^31-1)
--ως (2^31-1). Το εύρος τιμών μπορεί να αλλάξει με την χρήση της λέξης RANGE. Παράδειγμα
--ορισμού ενός σήματος με ακέραιη τιμή είναι το εξής:
signal m : integer range -32 to 32;
--Μια μεταβλητή τύπου integer με αρχική τιμή 0 και με όρια τιμών -128 έως 128 δηλώνεται ως εξής:
variable count : integer range -128 to 128 :=0;

--NATURAL Είναι υποτύπος του integer και περιλαμβάνει μη αρνητικούς ακεραίους (από 0 μέχρι
--και το άνω όριο των ακεραίων). Υποστηρίζει τις ίδιες πράξεις με τον τύπο integer.
--Παράδειγμα δήλωσης σήματος τύπου natural:
signal f : natural range 0 to 15;

--POSITIVE Είναι υποτύπος του integer και περιλαμβάνει μόνον θετικούς ακεραίους.

--BOOLEAN Ένα σήμα αυτού του τύπου μπορεί να πάρει την τιμή TRUE ή FALSE. Είναι
--βαθμωτός τύπος και υποστηρίζει λογικούς και σχεσιακούς τελεστές.

--CHARACTER Σήματα αυτού του τύπου μπορούν να πάρουν τιμές από ένα σύνολο 256
--συμβόλων των 8-bit. Τα σύμβολα αντιπροσωπεύουν το σύνολο χαρακτήρων ISO 8859-1, ενώ
--τα πρώτα 128 σύμβολα ανήκουν στον κοινό κώδικα ASCII. Αν και κάθε χαρακτήρας έχει
--εύρος 8 bits, ο τύπος διαχειρίζεται κάθε φορά ένα χαρακτήρα, οπότε είναι βαθμωτός.
--Υποστηρίζει σχεσιακούς τελεστές. Ο παράγωγος τύπος STRING ορίζεται ως πίνακας
--χαρακτήρων και υποστηρίζει σχεσιακούς τελεστές και τη συνένωση (concatenation ‘&’).

--TIME Αυτός ο τύπος δεδομένων προορίζεται μόνο για προσομοίωση (όχι για σύνθεση). Με τη
--βοήθειά του ορίζονται ακέραιοι, που παριστάνουν χρονικές στιγμές στον χρόνο προσομοίωσης.
--Υποστηρίζει τους αριθμητικούς και σχεσιακούς τελεστές.
