--Η αρχιτεκτονική (architecture) περιέχει µια ακριβή περιγραφή του τρόπου λειτουργίας του
--κυκλώµατος. Ξεκινά µε µια δήλωση: 

ARCHITECTURE όνοµα_αρχιτεκτονικής OF όνοµα_οντότητας IS 

--όπου όνοµα_αρχιτεκτονικής είναι ένα αλφαριθµητικό αναγνωριστικό, που ορίζει ο
--χρήστης για την αρχιτεκτονική και όνοµα_οντότητας είναι το ίδιο αναγνωριστικό µε το
--οποίο ο σχεδιαστής έχει ονοµάσει την οντότητα

--Η περιγραφή της αρχιτεκτονικής αρχίζει πάντα µε τη δεσµευµένη λέξη BEGIN. Τα σήµατα που
--ορίζονται στην οντότητα κληρονοµούνται στο σώµα της αρχιτεκτονικής µαζί µε τους τύπους
--τους. Ανάµεσα στη δήλωση της αρχιτεκτονικής και στη λέξη BEGIN µπορεί να υπάρχουν
--επιπλέον δηλώσεις σηµάτων εκτός από αυτά που έχουν δηλωθεί ως σήµατα εισόδων/εξόδων, τα
--οποία χρειάζονται για την περιγραφή της αρχιτεκτονικής.
--Άρα, η αρχιτεκτονική ενός κυκλώµατος σε VHDL περιγράφεται ως εξής: 

ARCHITECTURE όνοµα_αρχιτεκτονικής OF όνοµα_οντότητας IS
--[∆ηλώσεις επιπλέον σηµάτων]
BEGIN
--Εντολές που περιγράφουν λογικές λειτουργίες και αναθέτουν τιµές σε σήµατα
END [ARCHITECTURE] [όνοµα_αρχιτεκτονικής];
