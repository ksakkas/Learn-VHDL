--Χαρακτηριστικά (attributes)
--Η VHDL αποδίδει στους τύπους δεδομένων και στα αντικείμενα δεδομένων ορισμένα
--χαρακτηριστικά. Ένα χαρακτηριστικό μπορεί να είναι το κάτω ή το πάνω όριο της περιοχής ενός
--ακεραίου τύπου, ή η περιοχή δεικτών ενός τύπου πίνακα.
--(Διακρίνουμε χαρακτηριστικά βαθμωτών τύπων, χαρακτηριστικά τύπων πινάκων και
--χαρακτηριστικά σημάτων.

--Χαρακτηριστικά βαθμωτών τύπων
--Οι ακέραιοι τύποι είναι βαθμωτοί. Έστω ότι ένα τύπος integer έχει δηλωθεί ως εξής:
TYPE temp IS RANGE 0 to 273;
--Τότε, ορίζονται διάφορα χαρακτηριστικά του τύπου temp, που αναφέρονται ως:
<όνομα_τύπου>'<όνομα_χαρακτηριστικού> --, όπου η απόστροφος διαβάζεται “τικ”.
--Για παράδειγμα, το κάτω όριο της περιοχής τιμών του τύπου temp αναφέρεται ως temp'LOW
--και η τιμή του βέβαια είναι μηδέν. Η έκφραση:
Result<=temp'LOW --αναθέτει στο σήμα result την τιμή 0. Ο τύπος του σήματος result
--πρέπει να είναι temp.
--Αντίστοιχα, η έκφραση:
result<=temp'HIGH --, αναθέτει στο σήμα result την τιμή 273.
Το χαρακτηριστικό Temp'ASCENDING επιστρέφει TRUE αν η περιοχή τιμών του τύπου temp
είναι αύξουσα.

--Χαρακτηριστικά τύπων πίνακα (array)
--Έστω, τώρα, ότι έχει δηλωθεί από τον χρήστη ένας τύπος array δύο διαστάσεων, ως εξής:
TYPE TwoD IS ARRAY(0 to 10, 5 downto 0) OF std_logic_vector(3 downto 0);
--Μπορούν να αναζητηθούν οι τιμές χαρακτηριστικών του τύπου TwoD, όπως:
TwoD'LEFT(N) --, που σημαίνει «αριστερό όριο της νιοστής περιοχής δεικτών του τύπου πίνακα
--TwoD. Αν Ν=2, τότε η έκφραση y<= TwoD'LEFT(2) επιστρέφει στο σήμα y την τιμή 5. Το
--σήμα y πρέπει να είναι ίδιου τύπου όπως και η περιοχή τιμών, δηλαδή integer.

--Αντίστοιχα ορίζονται τα χαρακτηριστικά TwoD'RIGHT(N), TwoD'LOW(N) κι έχουν ακέραιη
--τιμή 10 και 0 αντίστοιχα, για Ν=1. Το χαρακτηριστικό TwoD'HIGH(2) έχει τιμή 5. Ας
--σημειωθεί ότι σε μονοδιάστατο πίνακα η παρένθεση (Ν) μπορεί να παραληφθεί.
--Τα παραπάνω χαρακτηριστικά μπορούν να πάρουν μέρος σε γενικευμένες δομές επανάληψης,
--όπως
FOR i IN x'LEFT to x'RIGHT LOOP…
--Εναλλακτικά, η παραπάνω επαναληπτική δομή μπορεί να γραφεί με τη βοήθεια του
--χαρακτηριστικού x'RANGE ως εξής:
FOR i IN x'RANGE LOOP…

--Χαρακτηριστικά σημάτων
--Το βασικότερο χαρακτηριστικό των σημάτων και αυτό που κυρίως χρησιμοποιούμε
--είναι το 'EVENT. Σημαίνει τη μετάβαση του σήματος και λαμβάνει τιμές TRUE ή FALSE:
SIGNAL s : std_logic;

--To χαρακτηριστικό s'EVENT λαμβάνει την τιμή TRUE αν κατά τη διάρκεια του παρόντος
--κύκλου έγινε μετάβαση του σήματος s από μια κατάσταση σε άλλη (π.χ. από '0' σε '1').
--Χρησιμοποιείται κατά κόρο σε ακολουθιακά συστήματα για να σημάνει τη μετάβαση σημάτων
--ρολογιού. Για παράδειγμα, έστω ότι σε ένα flip-flop έχει οριστεί σήμα clk τύπου std_logic.
--Τότε, η διατύπωση
IF clk'EVENT AND clk='1' THEN

--σημαίνει ότι η συνθήκη της IF αληθεύει αν έχει συμβεί μετάβαση ρολογιού
--(clk'EVENT=TRUE) ΚΑΙ η μετάβαση αυτή είναι απο το '0' στο '1'. Με άλλα λόγια η
--συνθήκη αληθεύει σε κάθε θετικό μέτωπο του παλμού ρολογιού.

